library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom_palette is
    generic(
        ADDR_WIDTH   : integer := 8
    );
    port (
        clk  : in std_logic;
        addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
        data : out std_logic_vector(23 downto 0)
    );
end rom_palette;

architecture rtl of rom_palette is
    type rom256x8 is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(23 downto 0); 
    constant romData : rom256x8 := (
         x"000000",
			x"002D00",
			x"003C00",
			x"006800",
			x"009800",
			x"00C400",
			x"00D300",
			x"00FF00",
			x"2D0000",
			x"2D2D00",
			x"2D3C00",
			x"2D6800",
			x"2D9800",
			x"2DC400",
			x"2DD300",
			x"2DFF00",
			x"470000",
			x"472D00",
			x"473C00",
			x"476800",
			x"479800",
			x"47C400",
			x"47D300",
			x"47FF00",
			x"730000",
			x"732D00",
			x"733C00",
			x"736800",
			x"739800",
			x"73C400",
			x"73D300",
			x"73FF00",
			x"8D0000",
			x"8D2D00",
			x"8D3C00",
			x"8D6800",
			x"8D9800",
			x"8DC400",
			x"8DD300",
			x"8DFF00",
			x"B90000",
			x"B92D00",
			x"B93C00",
			x"B96800",
			x"B99800",
			x"B9C400",
			x"B9D300",
			x"B9FF00",
			x"D30000",
			x"D32D00",
			x"D33C00",
			x"D36800",
			x"D39800",
			x"D3C400",
			x"D3D300",
			x"D3FF00",
			x"FF0000",
			x"FF2D00",
			x"FF3C00",
			x"FF6800",
			x"FF9800",
			x"FFC400",
			x"FFD300",
			x"FFFF00",
			x"00005B",
			x"002D5B",
			x"003C5B",
			x"00685B",
			x"00985B",
			x"00C45B",
			x"00D35B",
			x"00FF5B",
			x"2D005B",
			x"2D2D5B",
			x"2D3C5B",
			x"2D685B",
			x"2D985B",
			x"2DC45B",
			x"2DD35B",
			x"2DFF5B",
			x"47005B",
			x"472D5B",
			x"473C5B",
			x"47685B",
			x"47985B",
			x"47C45B",
			x"47D35B",
			x"47FF5B",
			x"73005B",
			x"732D5B",
			x"733C5B",
			x"73685B",
			x"73985B",
			x"73C45B",
			x"73D35B",
			x"73FF5B",
			x"8D005B",
			x"8D2D5B",
			x"8D3C5B",
			x"8D685B",
			x"8D985B",
			x"8DC45B",
			x"8DD35B",
			x"8DFF5B",
			x"B9005B",
			x"B92D5B",
			x"B93C5B",
			x"B9685B",
			x"B9985B",
			x"B9C45B",
			x"B9D35B",
			x"B9FF5B",
			x"D3005B",
			x"D32D5B",
			x"D33C5B",
			x"D3685B",
			x"D3985B",
			x"D3C45B",
			x"D3D35B",
			x"D3FF5B",
			x"FF005B",
			x"FF2D5B",
			x"FF3C5B",
			x"FF685B",
			x"FF985B",
			x"FFC45B",
			x"FFD35B",
			x"FFFF5B",
			x"0000A5",
			x"002DA5",
			x"003CA5",
			x"0068A5",
			x"0098A5",
			x"00C4A5",
			x"00D3A5",
			x"00FFA5",
			x"2D00A5",
			x"2D2DA5",
			x"2D3CA5",
			x"2D68A5",
			x"2D98A5",
			x"2DC4A5",
			x"2DD3A5",
			x"2DFFA5",
			x"4700A5",
			x"472DA5",
			x"473CA5",
			x"4768A5",
			x"4798A5",
			x"47C4A5",
			x"47D3A5",
			x"47FFA5",
			x"7300A5",
			x"732DA5",
			x"733CA5",
			x"7368A5",
			x"7398A5",
			x"73C4A5",
			x"73D3A5",
			x"73FFA5",
			x"8D00A5",
			x"8D2DA5",
			x"8D3CA5",
			x"8D68A5",
			x"8D98A5",
			x"8DC4A5",
			x"8DD3A5",
			x"8DFFA5",
			x"B900A5",
			x"B92DA5",
			x"B93CA5",
			x"B968A5",
			x"B998A5",
			x"B9C4A5",
			x"B9D3A5",
			x"B9FFA5",
			x"D300A5",
			x"D32DA5",
			x"D33CA5",
			x"D368A5",
			x"D398A5",
			x"D3C4A5",
			x"D3D3A5",
			x"D3FFA5",
			x"FF00A5",
			x"FF2DA5",
			x"FF3CA5",
			x"FF68A5",
			x"FF98A5",
			x"FFC4A5",
			x"FFD3A5",
			x"FFFFA5",
			x"0000FF",
			x"002DFF",
			x"003CFF",
			x"0068FF",
			x"0098FF",
			x"00C4FF",
			x"00D3FF",
			x"00FFFF",
			x"2D00FF",
			x"2D2DFF",
			x"2D3CFF",
			x"2D68FF",
			x"2D98FF",
			x"2DC4FF",
			x"2DD3FF",
			x"2DFFFF",
			x"4700FF",
			x"472DFF",
			x"473CFF",
			x"4768FF",
			x"4798FF",
			x"47C4FF",
			x"47D3FF",
			x"47FFFF",
			x"7300FF",
			x"732DFF",
			x"733CFF",
			x"7368FF",
			x"7398FF",
			x"73C4FF",
			x"73D3FF",
			x"73FFFF",
			x"8D00FF",
			x"8D2DFF",
			x"8D3CFF",
			x"8D68FF",
			x"8D98FF",
			x"8DC4FF",
			x"8DD3FF",
			x"8DFFFF",
			x"B900FF",
			x"B92DFF",
			x"B93CFF",
			x"B968FF",
			x"B998FF",
			x"B9C4FF",
			x"B9D3FF",
			x"B9FFFF",
			x"D300FF",
			x"D32DFF",
			x"D33CFF",
			x"D368FF",
			x"D398FF",
			x"D3C4FF",
			x"D3D3FF",
			x"D3FFFF",
			x"FF00FF",
			x"FF2DFF",
			x"FF3CFF",
			x"FF68FF",
			x"FF98FF",
			x"FFC4FF",
			x"FFD3FF",
			x"FFFFFF"
        );
    
begin
    process begin
        wait until rising_edge(clk);
        data <= romData(to_integer(unsigned(addr)));
    end process;
end;
